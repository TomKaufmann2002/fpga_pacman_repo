package font_pkg;

localparam [0:255][0:15][0:7] FONT = '{
    //   0 ' '
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //   1 '☺'
    '{
      8'b00000000,
      8'b00000000,
      8'b01111110,
      8'b10000001,
      8'b10100101,
      8'b10000001,
      8'b10000001,
      8'b10111101,
      8'b10011001,
      8'b10000001,
      8'b10000001,
      8'b01111110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //   2 '☻'
    '{
      8'b00000000,
      8'b00000000,
      8'b01111110,
      8'b11111111,
      8'b11011011,
      8'b11111111,
      8'b11111111,
      8'b11000011,
      8'b11100111,
      8'b11111111,
      8'b11111111,
      8'b01111110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //   3 '♥'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b01101100,
      8'b11111110,
      8'b11111110,
      8'b11111110,
      8'b11111110,
      8'b01111100,
      8'b00111000,
      8'b00010000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //   4 '♦'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00010000,
      8'b00111000,
      8'b01111100,
      8'b11111110,
      8'b01111100,
      8'b00111000,
      8'b00010000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //   5 '♣'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00011000,
      8'b00111100,
      8'b00111100,
      8'b11100111,
      8'b11100111,
      8'b11100111,
      8'b00011000,
      8'b00011000,
      8'b00111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //   6 '♠'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00011000,
      8'b00111100,
      8'b01111110,
      8'b11111111,
      8'b11111111,
      8'b01111110,
      8'b00011000,
      8'b00011000,
      8'b00111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //   7 '•'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00011000,
      8'b00111100,
      8'b00111100,
      8'b00011000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //   8 '◘'
    '{
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11100111,
      8'b11000011,
      8'b11000011,
      8'b11100111,
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11111111
    },
    //   9 '○'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00111100,
      8'b01100110,
      8'b01000010,
      8'b01000010,
      8'b01100110,
      8'b00111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  10 '◙'
    '{
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11000011,
      8'b10011001,
      8'b10111101,
      8'b10111101,
      8'b10011001,
      8'b11000011,
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11111111
    },
    //  11 '♂'
    '{
      8'b00000000,
      8'b00000000,
      8'b00011110,
      8'b00001110,
      8'b00011010,
      8'b00110010,
      8'b01111000,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b01111000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  12 '♀'
    '{
      8'b00000000,
      8'b00000000,
      8'b00111100,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b00111100,
      8'b00011000,
      8'b01111110,
      8'b00011000,
      8'b00011000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  13 '♪'
    '{
      8'b00000000,
      8'b00000000,
      8'b00111111,
      8'b00110011,
      8'b00111111,
      8'b00110000,
      8'b00110000,
      8'b00110000,
      8'b00110000,
      8'b01110000,
      8'b11110000,
      8'b11100000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  14 '♫'
    '{
      8'b00000000,
      8'b00000000,
      8'b01111111,
      8'b01100011,
      8'b01111111,
      8'b01100011,
      8'b01100011,
      8'b01100011,
      8'b01100011,
      8'b01100111,
      8'b11100111,
      8'b11100110,
      8'b11000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  15 '☼'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00011000,
      8'b00011000,
      8'b11011011,
      8'b00111100,
      8'b11100111,
      8'b00111100,
      8'b11011011,
      8'b00011000,
      8'b00011000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  16 '►'
    '{
      8'b00000000,
      8'b10000000,
      8'b11000000,
      8'b11100000,
      8'b11110000,
      8'b11111000,
      8'b11111110,
      8'b11111000,
      8'b11110000,
      8'b11100000,
      8'b11000000,
      8'b10000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  17 '◄'
    '{
      8'b00000000,
      8'b00000010,
      8'b00000110,
      8'b00001110,
      8'b00011110,
      8'b00111110,
      8'b11111110,
      8'b00111110,
      8'b00011110,
      8'b00001110,
      8'b00000110,
      8'b00000010,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  18 '↕'
    '{
      8'b00000000,
      8'b00000000,
      8'b00011000,
      8'b00111100,
      8'b01111110,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b01111110,
      8'b00111100,
      8'b00011000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  19 '‼'
    '{
      8'b00000000,
      8'b00000000,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b00000000,
      8'b01100110,
      8'b01100110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  20 '¶'
    '{
      8'b00000000,
      8'b00000000,
      8'b01111111,
      8'b11011011,
      8'b11011011,
      8'b11011011,
      8'b01111011,
      8'b00011011,
      8'b00011011,
      8'b00011011,
      8'b00011011,
      8'b00011011,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  21 '§'
    '{
      8'b00000000,
      8'b01111100,
      8'b11000110,
      8'b01100000,
      8'b00111000,
      8'b01101100,
      8'b11000110,
      8'b11000110,
      8'b01101100,
      8'b00111000,
      8'b00001100,
      8'b11000110,
      8'b01111100,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  22 '▬'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b11111110,
      8'b11111110,
      8'b11111110,
      8'b11111110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  23 '↨'
    '{
      8'b00000000,
      8'b00000000,
      8'b00011000,
      8'b00111100,
      8'b01111110,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b01111110,
      8'b00111100,
      8'b00011000,
      8'b01111110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  24 '↑'
    '{
      8'b00000000,
      8'b00000000,
      8'b00011000,
      8'b00111100,
      8'b01111110,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  25 '↓'
    '{
      8'b00000000,
      8'b00000000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b01111110,
      8'b00111100,
      8'b00011000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  26 '→'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00011000,
      8'b00001100,
      8'b11111110,
      8'b00001100,
      8'b00011000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  27 '←'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00110000,
      8'b01100000,
      8'b11111110,
      8'b01100000,
      8'b00110000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  28 '∟'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b11000000,
      8'b11000000,
      8'b11000000,
      8'b11111110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  29 '↔'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00101000,
      8'b01101100,
      8'b11111110,
      8'b01101100,
      8'b00101000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  30 '▲'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00010000,
      8'b00111000,
      8'b00111000,
      8'b01111100,
      8'b01111100,
      8'b11111110,
      8'b11111110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  31 '▼'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b11111110,
      8'b11111110,
      8'b01111100,
      8'b01111100,
      8'b00111000,
      8'b00111000,
      8'b00010000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  32 ' '
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  33 '!'
    '{
      8'b00000000,
      8'b00000000,
      8'b00011000,
      8'b00111100,
      8'b00111100,
      8'b00111100,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00000000,
      8'b00011000,
      8'b00011000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  34 '"'
    '{
      8'b00000000,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b00100100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  35 '#'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b01101100,
      8'b01101100,
      8'b11111110,
      8'b01101100,
      8'b01101100,
      8'b01101100,
      8'b11111110,
      8'b01101100,
      8'b01101100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  36 '$'
    '{
      8'b00011000,
      8'b00011000,
      8'b01111100,
      8'b11000110,
      8'b11000010,
      8'b11000000,
      8'b01111100,
      8'b00000110,
      8'b00000110,
      8'b10000110,
      8'b11000110,
      8'b01111100,
      8'b00011000,
      8'b00011000,
      8'b00000000,
      8'b00000000
    },
    //  37 '%'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b11000010,
      8'b11000110,
      8'b00001100,
      8'b00011000,
      8'b00110000,
      8'b01100000,
      8'b11000110,
      8'b10000110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  38 '&'
    '{
      8'b00000000,
      8'b00000000,
      8'b00111000,
      8'b01101100,
      8'b01101100,
      8'b00111000,
      8'b01110110,
      8'b11011100,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b01110110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  39 '\''
    '{
      8'b00000000,
      8'b00110000,
      8'b00110000,
      8'b00110000,
      8'b01100000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  40 '('
    '{
      8'b00000000,
      8'b00000000,
      8'b00001100,
      8'b00011000,
      8'b00110000,
      8'b00110000,
      8'b00110000,
      8'b00110000,
      8'b00110000,
      8'b00110000,
      8'b00011000,
      8'b00001100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  41 ')'
    '{
      8'b00000000,
      8'b00000000,
      8'b00110000,
      8'b00011000,
      8'b00001100,
      8'b00001100,
      8'b00001100,
      8'b00001100,
      8'b00001100,
      8'b00001100,
      8'b00011000,
      8'b00110000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  42 '*'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b01100110,
      8'b00111100,
      8'b11111111,
      8'b00111100,
      8'b01100110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  43 '+'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00011000,
      8'b00011000,
      8'b01111110,
      8'b00011000,
      8'b00011000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  44 ','
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00110000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  45 '-'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b11111110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  46 '.'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00011000,
      8'b00011000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  47 '/'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000010,
      8'b00000110,
      8'b00001100,
      8'b00011000,
      8'b00110000,
      8'b01100000,
      8'b11000000,
      8'b10000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  48 '0'
    '{
      8'b00000000,
      8'b00000000,
      8'b00111000,
      8'b01101100,
      8'b11000110,
      8'b11000110,
      8'b11010110,
      8'b11010110,
      8'b11000110,
      8'b11000110,
      8'b01101100,
      8'b00111000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  49 '1'
    '{
      8'b00000000,
      8'b00000000,
      8'b00011000,
      8'b00111000,
      8'b01111000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b01111110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  50 '2'
    '{
      8'b00000000,
      8'b00000000,
      8'b01111100,
      8'b11000110,
      8'b00000110,
      8'b00001100,
      8'b00011000,
      8'b00110000,
      8'b01100000,
      8'b11000000,
      8'b11000110,
      8'b11111110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  51 '3'
    '{
      8'b00000000,
      8'b00000000,
      8'b01111100,
      8'b11000110,
      8'b00000110,
      8'b00000110,
      8'b00111100,
      8'b00000110,
      8'b00000110,
      8'b00000110,
      8'b11000110,
      8'b01111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  52 '4'
    '{
      8'b00000000,
      8'b00000000,
      8'b00001100,
      8'b00011100,
      8'b00111100,
      8'b01101100,
      8'b11001100,
      8'b11111110,
      8'b00001100,
      8'b00001100,
      8'b00001100,
      8'b00011110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  53 '5'
    '{
      8'b00000000,
      8'b00000000,
      8'b11111110,
      8'b11000000,
      8'b11000000,
      8'b11000000,
      8'b11111100,
      8'b00000110,
      8'b00000110,
      8'b00000110,
      8'b11000110,
      8'b01111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  54 '6'
    '{
      8'b00000000,
      8'b00000000,
      8'b00111000,
      8'b01100000,
      8'b11000000,
      8'b11000000,
      8'b11111100,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b01111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  55 '7'
    '{
      8'b00000000,
      8'b00000000,
      8'b11111110,
      8'b11000110,
      8'b00000110,
      8'b00000110,
      8'b00001100,
      8'b00011000,
      8'b00110000,
      8'b00110000,
      8'b00110000,
      8'b00110000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  56 '8'
    '{
      8'b00000000,
      8'b00000000,
      8'b01111100,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b01111100,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b01111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  57 '9'
    '{
      8'b00000000,
      8'b00000000,
      8'b01111100,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b01111110,
      8'b00000110,
      8'b00000110,
      8'b00000110,
      8'b00001100,
      8'b01111000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  58 ':'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00011000,
      8'b00011000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00011000,
      8'b00011000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  59 ';'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00011000,
      8'b00011000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00011000,
      8'b00011000,
      8'b00110000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  60 '<'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000110,
      8'b00001100,
      8'b00011000,
      8'b00110000,
      8'b01100000,
      8'b00110000,
      8'b00011000,
      8'b00001100,
      8'b00000110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  61 '='
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b01111110,
      8'b00000000,
      8'b00000000,
      8'b01111110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  62 '>'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b01100000,
      8'b00110000,
      8'b00011000,
      8'b00001100,
      8'b00000110,
      8'b00001100,
      8'b00011000,
      8'b00110000,
      8'b01100000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  63 '?'
    '{
      8'b00000000,
      8'b00000000,
      8'b01111100,
      8'b11000110,
      8'b11000110,
      8'b00001100,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00000000,
      8'b00011000,
      8'b00011000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  64 '@'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b01111100,
      8'b11000110,
      8'b11000110,
      8'b11011110,
      8'b11011110,
      8'b11011110,
      8'b11011100,
      8'b11000000,
      8'b01111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  65 'A'
    '{
      8'b00000000,
      8'b00000000,
      8'b00010000,
      8'b00111000,
      8'b01101100,
      8'b11000110,
      8'b11000110,
      8'b11111110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  66 'B'
    '{
      8'b00000000,
      8'b00000000,
      8'b11111100,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b01111100,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b11111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  67 'C'
    '{
      8'b00000000,
      8'b00000000,
      8'b00111100,
      8'b01100110,
      8'b11000010,
      8'b11000000,
      8'b11000000,
      8'b11000000,
      8'b11000000,
      8'b11000010,
      8'b01100110,
      8'b00111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  68 'D'
    '{
      8'b00000000,
      8'b00000000,
      8'b11111000,
      8'b01101100,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b01101100,
      8'b11111000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  69 'E'
    '{
      8'b00000000,
      8'b00000000,
      8'b11111110,
      8'b01100110,
      8'b01100010,
      8'b01101000,
      8'b01111000,
      8'b01101000,
      8'b01100000,
      8'b01100010,
      8'b01100110,
      8'b11111110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  70 'F'
    '{
      8'b00000000,
      8'b00000000,
      8'b11111110,
      8'b01100110,
      8'b01100010,
      8'b01101000,
      8'b01111000,
      8'b01101000,
      8'b01100000,
      8'b01100000,
      8'b01100000,
      8'b11110000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  71 'G'
    '{
      8'b00000000,
      8'b00000000,
      8'b00111100,
      8'b01100110,
      8'b11000010,
      8'b11000000,
      8'b11000000,
      8'b11011110,
      8'b11000110,
      8'b11000110,
      8'b01100110,
      8'b00111010,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  72 'H'
    '{
      8'b00000000,
      8'b00000000,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11111110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  73 'I'
    '{
      8'b00000000,
      8'b00000000,
      8'b00111100,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  74 'J'
    '{
      8'b00000000,
      8'b00000000,
      8'b00011110,
      8'b00001100,
      8'b00001100,
      8'b00001100,
      8'b00001100,
      8'b00001100,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b01111000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  75 'K'
    '{
      8'b00000000,
      8'b00000000,
      8'b11100110,
      8'b01100110,
      8'b01100110,
      8'b01101100,
      8'b01111000,
      8'b01111000,
      8'b01101100,
      8'b01100110,
      8'b01100110,
      8'b11100110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  76 'L'
    '{
      8'b00000000,
      8'b00000000,
      8'b11110000,
      8'b01100000,
      8'b01100000,
      8'b01100000,
      8'b01100000,
      8'b01100000,
      8'b01100000,
      8'b01100010,
      8'b01100110,
      8'b11111110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  77 'M'
    '{
      8'b00000000,
      8'b00000000,
      8'b11000110,
      8'b11101110,
      8'b11111110,
      8'b11111110,
      8'b11010110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  78 'N'
    '{
      8'b00000000,
      8'b00000000,
      8'b11000110,
      8'b11100110,
      8'b11110110,
      8'b11111110,
      8'b11011110,
      8'b11001110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  79 'O'
    '{
      8'b00000000,
      8'b00000000,
      8'b01111100,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b01111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  80 'P'
    '{
      8'b00000000,
      8'b00000000,
      8'b11111100,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b01111100,
      8'b01100000,
      8'b01100000,
      8'b01100000,
      8'b01100000,
      8'b11110000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  81 'Q'
    '{
      8'b00000000,
      8'b00000000,
      8'b01111100,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11010110,
      8'b11011110,
      8'b01111100,
      8'b00001100,
      8'b00001110,
      8'b00000000,
      8'b00000000
    },
    //  82 'R'
    '{
      8'b00000000,
      8'b00000000,
      8'b11111100,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b01111100,
      8'b01101100,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b11100110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  83 'S'
    '{
      8'b00000000,
      8'b00000000,
      8'b01111100,
      8'b11000110,
      8'b11000110,
      8'b01100000,
      8'b00111000,
      8'b00001100,
      8'b00000110,
      8'b11000110,
      8'b11000110,
      8'b01111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  84 'T'
    '{
      8'b00000000,
      8'b00000000,
      8'b01111110,
      8'b01111110,
      8'b01011010,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  85 'U'
    '{
      8'b00000000,
      8'b00000000,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b01111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  86 'V'
    '{
      8'b00000000,
      8'b00000000,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b01101100,
      8'b00111000,
      8'b00010000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  87 'W'
    '{
      8'b00000000,
      8'b00000000,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11010110,
      8'b11010110,
      8'b11010110,
      8'b11111110,
      8'b11101110,
      8'b01101100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  88 'X'
    '{
      8'b00000000,
      8'b00000000,
      8'b11000110,
      8'b11000110,
      8'b01101100,
      8'b01111100,
      8'b00111000,
      8'b00111000,
      8'b01111100,
      8'b01101100,
      8'b11000110,
      8'b11000110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  89 'Y'
    '{
      8'b00000000,
      8'b00000000,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b00111100,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  90 'Z'
    '{
      8'b00000000,
      8'b00000000,
      8'b11111110,
      8'b11000110,
      8'b10000110,
      8'b00001100,
      8'b00011000,
      8'b00110000,
      8'b01100000,
      8'b11000010,
      8'b11000110,
      8'b11111110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  91 '['
    '{
      8'b00000000,
      8'b00000000,
      8'b00111100,
      8'b00110000,
      8'b00110000,
      8'b00110000,
      8'b00110000,
      8'b00110000,
      8'b00110000,
      8'b00110000,
      8'b00110000,
      8'b00111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  92 '\'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b10000000,
      8'b11000000,
      8'b11100000,
      8'b01110000,
      8'b00111000,
      8'b00011100,
      8'b00001110,
      8'b00000110,
      8'b00000010,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  93 ']'
    '{
      8'b00000000,
      8'b00000000,
      8'b00111100,
      8'b00001100,
      8'b00001100,
      8'b00001100,
      8'b00001100,
      8'b00001100,
      8'b00001100,
      8'b00001100,
      8'b00001100,
      8'b00111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  94 '^'
    '{
      8'b00010000,
      8'b00111000,
      8'b01101100,
      8'b11000110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  95 '_'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b11111111,
      8'b00000000,
      8'b00000000
    },
    //  96 '`'
    '{
      8'b00110000,
      8'b00110000,
      8'b00011000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  97 'a'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b01111000,
      8'b00001100,
      8'b01111100,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b01110110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  98 'b'
    '{
      8'b00000000,
      8'b00000000,
      8'b11100000,
      8'b01100000,
      8'b01100000,
      8'b01111000,
      8'b01101100,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b01111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    //  99 'c'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b01111100,
      8'b11000110,
      8'b11000000,
      8'b11000000,
      8'b11000000,
      8'b11000110,
      8'b01111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 100 'd'
    '{
      8'b00000000,
      8'b00000000,
      8'b00011100,
      8'b00001100,
      8'b00001100,
      8'b00111100,
      8'b01101100,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b01110110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 101 'e'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b01111100,
      8'b11000110,
      8'b11111110,
      8'b11000000,
      8'b11000000,
      8'b11000110,
      8'b01111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 102 'f'
    '{
      8'b00000000,
      8'b00000000,
      8'b00111000,
      8'b01101100,
      8'b01100100,
      8'b01100000,
      8'b11110000,
      8'b01100000,
      8'b01100000,
      8'b01100000,
      8'b01100000,
      8'b11110000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 103 'g'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b01110110,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b01111100,
      8'b00001100,
      8'b11001100,
      8'b01111000,
      8'b00000000
    },
    // 104 'h'
    '{
      8'b00000000,
      8'b00000000,
      8'b11100000,
      8'b01100000,
      8'b01100000,
      8'b01101100,
      8'b01110110,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b11100110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 105 'i'
    '{
      8'b00000000,
      8'b00000000,
      8'b00011000,
      8'b00011000,
      8'b00000000,
      8'b00111000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 106 'j'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000110,
      8'b00000110,
      8'b00000000,
      8'b00001110,
      8'b00000110,
      8'b00000110,
      8'b00000110,
      8'b00000110,
      8'b00000110,
      8'b00000110,
      8'b01100110,
      8'b01100110,
      8'b00111100,
      8'b00000000
    },
    // 107 'k'
    '{
      8'b00000000,
      8'b00000000,
      8'b11100000,
      8'b01100000,
      8'b01100000,
      8'b01100110,
      8'b01101100,
      8'b01111000,
      8'b01111000,
      8'b01101100,
      8'b01100110,
      8'b11100110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 108 'l'
    '{
      8'b00000000,
      8'b00000000,
      8'b00111000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 109 'm'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b11101100,
      8'b11111110,
      8'b11010110,
      8'b11010110,
      8'b11010110,
      8'b11010110,
      8'b11000110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 110 'n'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b11011100,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 111 'o'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b01111100,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b01111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 112 'p'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b11011100,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b01111100,
      8'b01100000,
      8'b01100000,
      8'b11110000,
      8'b00000000
    },
    // 113 'q'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b01110110,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b01111100,
      8'b00001100,
      8'b00001100,
      8'b00011110,
      8'b00000000
    },
    // 114 'r'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b11011100,
      8'b01110110,
      8'b01100110,
      8'b01100000,
      8'b01100000,
      8'b01100000,
      8'b11110000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 115 's'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b01111100,
      8'b11000110,
      8'b01100000,
      8'b00111000,
      8'b00001100,
      8'b11000110,
      8'b01111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 116 't'
    '{
      8'b00000000,
      8'b00000000,
      8'b00010000,
      8'b00110000,
      8'b00110000,
      8'b11111100,
      8'b00110000,
      8'b00110000,
      8'b00110000,
      8'b00110000,
      8'b00110110,
      8'b00011100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 117 'u'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b01110110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 118 'v'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b00111100,
      8'b00011000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 119 'w'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b11000110,
      8'b11000110,
      8'b11010110,
      8'b11010110,
      8'b11010110,
      8'b11111110,
      8'b01101100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 120 'x'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b11000110,
      8'b01101100,
      8'b00111000,
      8'b00111000,
      8'b00111000,
      8'b01101100,
      8'b11000110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 121 'y'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b01111110,
      8'b00000110,
      8'b00001100,
      8'b11111000,
      8'b00000000
    },
    // 122 'z'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b11111110,
      8'b11001100,
      8'b00011000,
      8'b00110000,
      8'b01100000,
      8'b11000110,
      8'b11111110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 123 '{'
    '{
      8'b00000000,
      8'b00000000,
      8'b00001110,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b01110000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00001110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 124 '|'
    '{
      8'b00000000,
      8'b00000000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00000000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 125 '}'
    '{
      8'b00000000,
      8'b00000000,
      8'b01110000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00001110,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b01110000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 126 '~'
    '{
      8'b00000000,
      8'b00000000,
      8'b01110110,
      8'b11011100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 127 '⌂'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00010000,
      8'b00111000,
      8'b01101100,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11111110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 128 'Ç'
    '{
      8'b00000000,
      8'b00000000,
      8'b00111100,
      8'b01100110,
      8'b11000010,
      8'b11000000,
      8'b11000000,
      8'b11000000,
      8'b11000010,
      8'b01100110,
      8'b00111100,
      8'b00001100,
      8'b00000110,
      8'b01111100,
      8'b00000000,
      8'b00000000
    },
    // 129 'ü'
    '{
      8'b00000000,
      8'b00000000,
      8'b11001100,
      8'b00000000,
      8'b00000000,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b01110110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 130 'é'
    '{
      8'b00000000,
      8'b00001100,
      8'b00011000,
      8'b00110000,
      8'b00000000,
      8'b01111100,
      8'b11000110,
      8'b11111110,
      8'b11000000,
      8'b11000000,
      8'b11000110,
      8'b01111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 131 'â'
    '{
      8'b00000000,
      8'b00010000,
      8'b00111000,
      8'b01101100,
      8'b00000000,
      8'b01111000,
      8'b00001100,
      8'b01111100,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b01110110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 132 'ä'
    '{
      8'b00000000,
      8'b00000000,
      8'b11001100,
      8'b00000000,
      8'b00000000,
      8'b01111000,
      8'b00001100,
      8'b01111100,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b01110110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 133 'à'
    '{
      8'b00000000,
      8'b01100000,
      8'b00110000,
      8'b00011000,
      8'b00000000,
      8'b01111000,
      8'b00001100,
      8'b01111100,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b01110110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 134 'å'
    '{
      8'b00000000,
      8'b00111000,
      8'b01101100,
      8'b00111000,
      8'b00000000,
      8'b01111000,
      8'b00001100,
      8'b01111100,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b01110110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 135 'ç'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00111100,
      8'b01100110,
      8'b01100000,
      8'b01100000,
      8'b01100110,
      8'b00111100,
      8'b00001100,
      8'b00000110,
      8'b00111100,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 136 'ê'
    '{
      8'b00000000,
      8'b00010000,
      8'b00111000,
      8'b01101100,
      8'b00000000,
      8'b01111100,
      8'b11000110,
      8'b11111110,
      8'b11000000,
      8'b11000000,
      8'b11000110,
      8'b01111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 137 'ë'
    '{
      8'b00000000,
      8'b00000000,
      8'b11000110,
      8'b00000000,
      8'b00000000,
      8'b01111100,
      8'b11000110,
      8'b11111110,
      8'b11000000,
      8'b11000000,
      8'b11000110,
      8'b01111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 138 'è'
    '{
      8'b00000000,
      8'b01100000,
      8'b00110000,
      8'b00011000,
      8'b00000000,
      8'b01111100,
      8'b11000110,
      8'b11111110,
      8'b11000000,
      8'b11000000,
      8'b11000110,
      8'b01111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 139 'ï'
    '{
      8'b00000000,
      8'b00000000,
      8'b01100110,
      8'b00000000,
      8'b00000000,
      8'b00111000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 140 'î'
    '{
      8'b00000000,
      8'b00011000,
      8'b00111100,
      8'b01100110,
      8'b00000000,
      8'b00111000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 141 'ì'
    '{
      8'b00000000,
      8'b01100000,
      8'b00110000,
      8'b00011000,
      8'b00000000,
      8'b00111000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 142 'Ä'
    '{
      8'b00000000,
      8'b11000110,
      8'b00000000,
      8'b00010000,
      8'b00111000,
      8'b01101100,
      8'b11000110,
      8'b11000110,
      8'b11111110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 143 'Å'
    '{
      8'b00111000,
      8'b01101100,
      8'b00111000,
      8'b00000000,
      8'b00111000,
      8'b01101100,
      8'b11000110,
      8'b11000110,
      8'b11111110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 144 'É'
    '{
      8'b00011000,
      8'b00110000,
      8'b01100000,
      8'b00000000,
      8'b11111110,
      8'b01100110,
      8'b01100000,
      8'b01111100,
      8'b01100000,
      8'b01100000,
      8'b01100110,
      8'b11111110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 145 'æ'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b11001100,
      8'b01110110,
      8'b00110110,
      8'b01111110,
      8'b11011000,
      8'b11011000,
      8'b01101110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 146 'Æ'
    '{
      8'b00000000,
      8'b00000000,
      8'b00111110,
      8'b01101100,
      8'b11001100,
      8'b11001100,
      8'b11111110,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b11001110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 147 'ô'
    '{
      8'b00000000,
      8'b00010000,
      8'b00111000,
      8'b01101100,
      8'b00000000,
      8'b01111100,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b01111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 148 'ö'
    '{
      8'b00000000,
      8'b00000000,
      8'b11000110,
      8'b00000000,
      8'b00000000,
      8'b01111100,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b01111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 149 'ò'
    '{
      8'b00000000,
      8'b01100000,
      8'b00110000,
      8'b00011000,
      8'b00000000,
      8'b01111100,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b01111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 150 'û'
    '{
      8'b00000000,
      8'b00110000,
      8'b01111000,
      8'b11001100,
      8'b00000000,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b01110110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 151 'ù'
    '{
      8'b00000000,
      8'b01100000,
      8'b00110000,
      8'b00011000,
      8'b00000000,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b01110110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 152 'ÿ'
    '{
      8'b00000000,
      8'b00000000,
      8'b11000110,
      8'b00000000,
      8'b00000000,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b01111110,
      8'b00000110,
      8'b00001100,
      8'b01111000,
      8'b00000000
    },
    // 153 'Ö'
    '{
      8'b00000000,
      8'b11000110,
      8'b00000000,
      8'b01111100,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b01111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 154 'Ü'
    '{
      8'b00000000,
      8'b11000110,
      8'b00000000,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b01111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 155 '¢'
    '{
      8'b00000000,
      8'b00011000,
      8'b00011000,
      8'b00111100,
      8'b01100110,
      8'b01100000,
      8'b01100000,
      8'b01100000,
      8'b01100110,
      8'b00111100,
      8'b00011000,
      8'b00011000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 156 '£'
    '{
      8'b00000000,
      8'b00111000,
      8'b01101100,
      8'b01100100,
      8'b01100000,
      8'b11110000,
      8'b01100000,
      8'b01100000,
      8'b01100000,
      8'b01100000,
      8'b11100110,
      8'b11111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 157 '¥'
    '{
      8'b00000000,
      8'b00000000,
      8'b01100110,
      8'b01100110,
      8'b00111100,
      8'b00011000,
      8'b01111110,
      8'b00011000,
      8'b01111110,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 158 '₧'
    '{
      8'b00000000,
      8'b11111000,
      8'b11001100,
      8'b11001100,
      8'b11111000,
      8'b11000100,
      8'b11001100,
      8'b11011110,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b11000110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 159 'ƒ'
    '{
      8'b00000000,
      8'b00001110,
      8'b00011011,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b01111110,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b11011000,
      8'b01110000,
      8'b00000000,
      8'b00000000
    },
    // 160 'á'
    '{
      8'b00000000,
      8'b00011000,
      8'b00110000,
      8'b01100000,
      8'b00000000,
      8'b01111000,
      8'b00001100,
      8'b01111100,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b01110110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 161 'í'
    '{
      8'b00000000,
      8'b00001100,
      8'b00011000,
      8'b00110000,
      8'b00000000,
      8'b00111000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 162 'ó'
    '{
      8'b00000000,
      8'b00011000,
      8'b00110000,
      8'b01100000,
      8'b00000000,
      8'b01111100,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b01111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 163 'ú'
    '{
      8'b00000000,
      8'b00011000,
      8'b00110000,
      8'b01100000,
      8'b00000000,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b01110110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 164 'ñ'
    '{
      8'b00000000,
      8'b00000000,
      8'b01110110,
      8'b11011100,
      8'b00000000,
      8'b11011100,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 165 'Ñ'
    '{
      8'b01110110,
      8'b11011100,
      8'b00000000,
      8'b11000110,
      8'b11100110,
      8'b11110110,
      8'b11111110,
      8'b11011110,
      8'b11001110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 166 'ª'
    '{
      8'b00000000,
      8'b00111100,
      8'b01101100,
      8'b01101100,
      8'b00111110,
      8'b00000000,
      8'b01111110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 167 'º'
    '{
      8'b00000000,
      8'b00111000,
      8'b01101100,
      8'b01101100,
      8'b00111000,
      8'b00000000,
      8'b01111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 168 '¿'
    '{
      8'b00000000,
      8'b00000000,
      8'b00110000,
      8'b00110000,
      8'b00000000,
      8'b00110000,
      8'b00110000,
      8'b01100000,
      8'b11000000,
      8'b11000110,
      8'b11000110,
      8'b01111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 169 '⌐'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b11111110,
      8'b11000000,
      8'b11000000,
      8'b11000000,
      8'b11000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 170 '¬'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b11111110,
      8'b00000110,
      8'b00000110,
      8'b00000110,
      8'b00000110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 171 '½'
    '{
      8'b00000000,
      8'b11000000,
      8'b11000000,
      8'b11000010,
      8'b11000110,
      8'b11001100,
      8'b00011000,
      8'b00110000,
      8'b01100000,
      8'b11011100,
      8'b10000110,
      8'b00001100,
      8'b00011000,
      8'b00111110,
      8'b00000000,
      8'b00000000
    },
    // 172 '¼'
    '{
      8'b00000000,
      8'b11000000,
      8'b11000000,
      8'b11000010,
      8'b11000110,
      8'b11001100,
      8'b00011000,
      8'b00110000,
      8'b01100110,
      8'b11001110,
      8'b10011110,
      8'b00111110,
      8'b00000110,
      8'b00000110,
      8'b00000000,
      8'b00000000
    },
    // 173 '¡'
    '{
      8'b00000000,
      8'b00000000,
      8'b00011000,
      8'b00011000,
      8'b00000000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00111100,
      8'b00111100,
      8'b00111100,
      8'b00011000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 174 '«'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00110110,
      8'b01101100,
      8'b11011000,
      8'b01101100,
      8'b00110110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 175 '»'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b11011000,
      8'b01101100,
      8'b00110110,
      8'b01101100,
      8'b11011000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 176 '░'
    '{
      8'b00010001,
      8'b01000100,
      8'b00010001,
      8'b01000100,
      8'b00010001,
      8'b01000100,
      8'b00010001,
      8'b01000100,
      8'b00010001,
      8'b01000100,
      8'b00010001,
      8'b01000100,
      8'b00010001,
      8'b01000100,
      8'b00010001,
      8'b01000100
    },
    // 177 '▒'
    '{
      8'b01010101,
      8'b10101010,
      8'b01010101,
      8'b10101010,
      8'b01010101,
      8'b10101010,
      8'b01010101,
      8'b10101010,
      8'b01010101,
      8'b10101010,
      8'b01010101,
      8'b10101010,
      8'b01010101,
      8'b10101010,
      8'b01010101,
      8'b10101010
    },
    // 178 '▓'
    '{
      8'b11011101,
      8'b01110111,
      8'b11011101,
      8'b01110111,
      8'b11011101,
      8'b01110111,
      8'b11011101,
      8'b01110111,
      8'b11011101,
      8'b01110111,
      8'b11011101,
      8'b01110111,
      8'b11011101,
      8'b01110111,
      8'b11011101,
      8'b01110111
    },
    // 179 '│'
    '{
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000
    },
    // 180 '┤'
    '{
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b11111000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000
    },
    // 181 '╡'
    '{
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b11111000,
      8'b00011000,
      8'b11111000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000
    },
    // 182 '╢'
    '{
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b11110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110
    },
    // 183 '╖'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b11111110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110
    },
    // 184 '╕'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b11111000,
      8'b00011000,
      8'b11111000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000
    },
    // 185 '╣'
    '{
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b11110110,
      8'b00000110,
      8'b11110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110
    },
    // 186 '║'
    '{
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110
    },
    // 187 '╗'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b11111110,
      8'b00000110,
      8'b11110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110
    },
    // 188 '╝'
    '{
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b11110110,
      8'b00000110,
      8'b11111110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 189 '╜'
    '{
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b11111110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 190 '╛'
    '{
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b11111000,
      8'b00011000,
      8'b11111000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 191 '┐'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b11111000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000
    },
    // 192 '└'
    '{
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011111,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 193 '┴'
    '{
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b11111111,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 194 '┬'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b11111111,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000
    },
    // 195 '├'
    '{
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011111,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000
    },
    // 196 '─'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b11111111,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 197 '┼'
    '{
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b11111111,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000
    },
    // 198 '╞'
    '{
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011111,
      8'b00011000,
      8'b00011111,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000
    },
    // 199 '╟'
    '{
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110111,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110
    },
    // 200 '╚'
    '{
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110111,
      8'b00110000,
      8'b00111111,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 201 '╔'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00111111,
      8'b00110000,
      8'b00110111,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110
    },
    // 202 '╩'
    '{
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b11110111,
      8'b00000000,
      8'b11111111,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 203 '╦'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b11111111,
      8'b00000000,
      8'b11110111,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110
    },
    // 204 '╠'
    '{
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110111,
      8'b00110000,
      8'b00110111,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110
    },
    // 205 '═'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b11111111,
      8'b00000000,
      8'b11111111,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 206 '╬'
    '{
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b11110111,
      8'b00000000,
      8'b11110111,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110
    },
    // 207 '╧'
    '{
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b11111111,
      8'b00000000,
      8'b11111111,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 208 '╨'
    '{
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b11111111,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 209 '╤'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b11111111,
      8'b00000000,
      8'b11111111,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000
    },
    // 210 '╥'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b11111111,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110
    },
    // 211 '╙'
    '{
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00111111,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 212 '╘'
    '{
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011111,
      8'b00011000,
      8'b00011111,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 213 '╒'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00011111,
      8'b00011000,
      8'b00011111,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000
    },
    // 214 '╓'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00111111,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110
    },
    // 215 '╫'
    '{
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b11111111,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110,
      8'b00110110
    },
    // 216 '╪'
    '{
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b11111111,
      8'b00011000,
      8'b11111111,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000
    },
    // 217 '┘'
    '{
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b11111000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 218 '┌'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00011111,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000
    },
    // 219 '█'
    '{
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11111111
    },
    // 220 '▄'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11111111
    },
    // 221 '▌'
    '{
      8'b11110000,
      8'b11110000,
      8'b11110000,
      8'b11110000,
      8'b11110000,
      8'b11110000,
      8'b11110000,
      8'b11110000,
      8'b11110000,
      8'b11110000,
      8'b11110000,
      8'b11110000,
      8'b11110000,
      8'b11110000,
      8'b11110000,
      8'b11110000
    },
    // 222 '▐'
    '{
      8'b00001111,
      8'b00001111,
      8'b00001111,
      8'b00001111,
      8'b00001111,
      8'b00001111,
      8'b00001111,
      8'b00001111,
      8'b00001111,
      8'b00001111,
      8'b00001111,
      8'b00001111,
      8'b00001111,
      8'b00001111,
      8'b00001111,
      8'b00001111
    },
    // 223 '▀'
    '{
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b11111111,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 224 'α'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b01110110,
      8'b11011100,
      8'b11011000,
      8'b11011000,
      8'b11011000,
      8'b11011100,
      8'b01110110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 225 'ß'
    '{
      8'b00000000,
      8'b00000000,
      8'b01111000,
      8'b11001100,
      8'b11001100,
      8'b11001100,
      8'b11011000,
      8'b11001100,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11001100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 226 'Γ'
    '{
      8'b00000000,
      8'b00000000,
      8'b11111110,
      8'b11000110,
      8'b11000110,
      8'b11000000,
      8'b11000000,
      8'b11000000,
      8'b11000000,
      8'b11000000,
      8'b11000000,
      8'b11000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 227 'π'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b11111110,
      8'b01101100,
      8'b01101100,
      8'b01101100,
      8'b01101100,
      8'b01101100,
      8'b01101100,
      8'b01101100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 228 'Σ'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b11111110,
      8'b11000110,
      8'b01100000,
      8'b00110000,
      8'b00011000,
      8'b00110000,
      8'b01100000,
      8'b11000110,
      8'b11111110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 229 'σ'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b01111110,
      8'b11011000,
      8'b11011000,
      8'b11011000,
      8'b11011000,
      8'b11011000,
      8'b01110000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 230 'µ'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b01111100,
      8'b01100000,
      8'b01100000,
      8'b11000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 231 'τ'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b01110110,
      8'b11011100,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 232 'Φ'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b01111110,
      8'b00011000,
      8'b00111100,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b00111100,
      8'b00011000,
      8'b01111110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 233 'Θ'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00111000,
      8'b01101100,
      8'b11000110,
      8'b11000110,
      8'b11111110,
      8'b11000110,
      8'b11000110,
      8'b01101100,
      8'b00111000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 234 'Ω'
    '{
      8'b00000000,
      8'b00000000,
      8'b00111000,
      8'b01101100,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b01101100,
      8'b01101100,
      8'b01101100,
      8'b01101100,
      8'b11101110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 235 'δ'
    '{
      8'b00000000,
      8'b00000000,
      8'b00011110,
      8'b00110000,
      8'b00011000,
      8'b00001100,
      8'b00111110,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b01100110,
      8'b00111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 236 '∞'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b01111110,
      8'b11011011,
      8'b11011011,
      8'b11011011,
      8'b01111110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 237 'φ'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000011,
      8'b00000110,
      8'b01111110,
      8'b11011011,
      8'b11011011,
      8'b11110011,
      8'b01111110,
      8'b01100000,
      8'b11000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 238 'ε'
    '{
      8'b00000000,
      8'b00000000,
      8'b00011100,
      8'b00110000,
      8'b01100000,
      8'b01100000,
      8'b01111100,
      8'b01100000,
      8'b01100000,
      8'b01100000,
      8'b00110000,
      8'b00011100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 239 '∩'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b01111100,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b11000110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 240 '≡'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b11111110,
      8'b00000000,
      8'b00000000,
      8'b11111110,
      8'b00000000,
      8'b00000000,
      8'b11111110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 241 '±'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00011000,
      8'b00011000,
      8'b01111110,
      8'b00011000,
      8'b00011000,
      8'b00000000,
      8'b00000000,
      8'b11111111,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 242 '≥'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00110000,
      8'b00011000,
      8'b00001100,
      8'b00000110,
      8'b00001100,
      8'b00011000,
      8'b00110000,
      8'b00000000,
      8'b01111110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 243 '≤'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00001100,
      8'b00011000,
      8'b00110000,
      8'b01100000,
      8'b00110000,
      8'b00011000,
      8'b00001100,
      8'b00000000,
      8'b01111110,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 244 '⌠'
    '{
      8'b00000000,
      8'b00000000,
      8'b00001110,
      8'b00011011,
      8'b00011011,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000
    },
    // 245 '⌡'
    '{
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b00011000,
      8'b11011000,
      8'b11011000,
      8'b11011000,
      8'b01110000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 246 '÷'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00011000,
      8'b00011000,
      8'b00000000,
      8'b01111110,
      8'b00000000,
      8'b00011000,
      8'b00011000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 247 '≈'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b01110110,
      8'b11011100,
      8'b00000000,
      8'b01110110,
      8'b11011100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 248 '°'
    '{
      8'b00000000,
      8'b00111000,
      8'b01101100,
      8'b01101100,
      8'b00111000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 249 '∙'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00011000,
      8'b00011000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 250 '·'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00011000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 251 '√'
    '{
      8'b00000000,
      8'b00001111,
      8'b00001100,
      8'b00001100,
      8'b00001100,
      8'b00001100,
      8'b00001100,
      8'b11101100,
      8'b01101100,
      8'b01101100,
      8'b00111100,
      8'b00011100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 252 'ⁿ'
    '{
      8'b00000000,
      8'b11011000,
      8'b01101100,
      8'b01101100,
      8'b01101100,
      8'b01101100,
      8'b01101100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 253 '²'
    '{
      8'b00000000,
      8'b01110000,
      8'b11011000,
      8'b00110000,
      8'b01100000,
      8'b11001000,
      8'b11111000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 254 '■'
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b01111100,
      8'b01111100,
      8'b01111100,
      8'b01111100,
      8'b01111100,
      8'b01111100,
      8'b01111100,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    },
    // 255 ' '
    '{
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000,
      8'b00000000
    }
  };
  


endpackage
